library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity VGA is port (

			clk  		: in std_logic;
			clk1hz  		: in std_logic;
			q0,q1,q3    : in integer range 0 to 9;
			q2    : in integer range 0 to 5;
			estado : in integer range 0 to 8;
			flag  		: in std_logic;
			flag_fim  		: in std_logic;
			sync_h    	: out std_logic;
			sync_v    	: out std_logic;
			corestovga   	: out std_logic_vector(7 downto 0)
			);
end VGA;

architecture hardware of VGA is
-------------------------DEFINI��O DAS MATRIZES-------------------------------------------	
type digito is array (0 to 97) of std_logic_vector (0 to 63);
type ponto is array (0 to 97) of std_logic_vector (0 to 63);

-------------------------CONTANTES ATRIBUIDAS AS MATRIZES----------------------------------
--ABAIXO AS MATRIZES REPRESENTENADO 0,1,2,3,4,5,6,7,8,9 e '.'

constant digito0 : digito := (
	"0000000000000000000000000011111111111100000000000000000000000000",
	"0000000000000000000000111111111111111111110000000000000000000000",
	"0000000000000000000011111111111111111111111100000000000000000000",
	"0000000000000000001111111111111111111111111111000000000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000001111111111111111111111111111111111000000000000000",
	"0000000000000111111111111111111111111111111111111100000000000000",
	"0000000000001111111111111111111111111111111111111111000000000000",
	"0000000000011111111111111111111111111111111111111111000000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111100000011111111111111111111111000000",
	"0000001111111111111111111110000000000111111111111111111111000000",
	"0000001111111111111111111100000000000011111111111111111111000000",
	"0000011111111111111111111000000000000001111111111111111111100000",
	"0000011111111111111111110000000000000000111111111111111111100000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111000000000000000000001111111111111111110000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000011111111111111111100",
	"0011111111111111111100000000000000000000000011111111111111111100",
	"0011111111111111111100000000000000000000000011111111111111111100",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0011111111111111111100000000000000000000000011111111111111111100",
	"0011111111111111111100000000000000000000000011111111111111111100",
	"0011111111111111111100000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111110000000000000000000000111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000011111111111111111110000000000000000111111111111111111100000",
	"0000011111111111111111111000000000000001111111111111111111100000",
	"0000011111111111111111111100000000000011111111111111111111000000",
	"0000001111111111111111111110000000000111111111111111111111000000",
	"0000001111111111111111111111100000011111111111111111111111000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000000001111111111111111111111111111111111111111100000000000",
	"0000000000000111111111111111111111111111111111111111000000000000",
	"0000000000000011111111111111111111111111111111111110000000000000",
	"0000000000000001111111111111111111111111111111111000000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000000001111111111111111111111111111000000000000000000",
	"0000000000000000000011111111111111111111111100000000000000000000",
	"0000000000000000000000111111111111111111110000000000000000000000",
	"0000000000000000000000000011111111111100000000000000000000000000");
	
	
constant digito1 : digito := (
		"0000000000000000000000000000111111111111111000000000000000000000",
		"0000000000000000000000000000111111111111111000000000000000000000",
		"0000000000000000000000000001111111111111111000000000000000000000",
		"0000000000000000000000000001111111111111111000000000000000000000",
		"0000000000000000000000000011111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000001111111111111111111000000000000000000000",
		"0000000000000000000000011111111111111111111000000000000000000000",
		"0000000000000000000000011111111111111111111000000000000000000000",
		"0000000000000000000000111111111111111111111000000000000000000000",
		"0000000000000000000001111111111111111111111000000000000000000000",
		"0000000000000000000011111111111111111111111000000000000000000000",
		"0000000000000000000111111111111111111111111000000000000000000000",
		"0000000000000000011111111111111111111111111000000000000000000000",
		"0000000000000000111111111111111111111111111000000000000000000000",
		"0000000000000001111111111111111111111111111000000000000000000000",
		"0000000000000111111111111111111111111111111000000000000000000000",
		"0000000000001111111111111111111111111111111000000000000000000000",
		"0000000000111111111111111111111111111111111000000000000000000000",
		"0000000001111111111111111111111111111111111000000000000000000000",
		"0000000111111111111111111111111111111111111000000000000000000000",
		"0000011111111111111111111111111111111111111000000000000000000000",
		"0011111111111111111111111111111111111111111000000000000000000000",
		"0111111111111111111111111111111111111111111000000000000000000000",
		"0111111111111111111111111111111111111111111000000000000000000000",
		"0111111111111111111111111111111111111111111000000000000000000000",
		"0111111111111111111111110111111111111111111000000000000000000000",
		"0111111111111111111111100111111111111111111000000000000000000000",
		"0111111111111111111111000111111111111111111000000000000000000000",
		"0111111111111111111110000111111111111111111000000000000000000000",
		"0111111111111111111100000111111111111111111000000000000000000000",
		"0111111111111111111000000111111111111111111000000000000000000000",
		"0111111111111111100000000111111111111111111000000000000000000000",
		"0111111111111111000000000111111111111111111000000000000000000000",
		"0111111111111100000000000111111111111111111000000000000000000000",
		"0111111111111000000000000111111111111111111000000000000000000000",
		"0111111111100000000000000111111111111111111000000000000000000000",
		"0111111110000000000000000111111111111111111000000000000000000000",
		"0111111000000000000000000111111111111111111000000000000000000000",
		"0111100000000000000000000111111111111111111000000000000000000000",
		"0100000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000111111111111111111000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000");
	
	
	
	constant digito2 : digito := (
	"0000000000000000000000000001111111111111000000000000000000000000",
	"0000000000000000000000011111111111111111111110000000000000000000",
	"0000000000000000000011111111111111111111111111110000000000000000",
	"0000000000000000001111111111111111111111111111111100000000000000",
	"0000000000000000111111111111111111111111111111111110000000000000",
	"0000000000000011111111111111111111111111111111111111100000000000",
	"0000000000000111111111111111111111111111111111111111110000000000",
	"0000000000001111111111111111111111111111111111111111111000000000",
	"0000000000011111111111111111111111111111111111111111111100000000",
	"0000000000111111111111111111111111111111111111111111111110000000",
	"0000000001111111111111111111111111111111111111111111111111000000",
	"0000000011111111111111111111111111111111111111111111111111100000",
	"0000000011111111111111111111111111111111111111111111111111100000",
	"0000000111111111111111111111111111111111111111111111111111110000",
	"0000000111111111111111111111111111111111111111111111111111110000",
	"0000001111111111111111111111111111111111111111111111111111111000",
	"0000001111111111111111111111110000000111111111111111111111111000",
	"0000011111111111111111111110000000000001111111111111111111111100",
	"0000011111111111111111111100000000000000111111111111111111111100",
	"0000011111111111111111111000000000000000011111111111111111111100",
	"0000111111111111111111110000000000000000001111111111111111111100",
	"0000111111111111111111110000000000000000000111111111111111111110",
	"0000111111111111111111100000000000000000000111111111111111111110",
	"0000111111111111111111100000000000000000000111111111111111111110",
	"0000111111111111111111100000000000000000000011111111111111111110",
	"0001111111111111111111100000000000000000000011111111111111111110",
	"0001111111111111111111000000000000000000000011111111111111111110",
	"0001111111111111111111000000000000000000000011111111111111111110",
	"0000011111111111111111000000000000000000000011111111111111111110",
	"0000000000000000111111000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111100",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000001111111111111111111000",
	"0000000000000000000000000000000000000000001111111111111111111000",
	"0000000000000000000000000000000000000000011111111111111111111000",
	"0000000000000000000000000000000000000000011111111111111111110000",
	"0000000000000000000000000000000000000000111111111111111111110000",
	"0000000000000000000000000000000000000001111111111111111111100000",
	"0000000000000000000000000000000000000011111111111111111111100000",
	"0000000000000000000000000000000000000111111111111111111111000000",
	"0000000000000000000000000000000000000111111111111111111111000000",
	"0000000000000000000000000000000000001111111111111111111110000000",
	"0000000000000000000000000000000000011111111111111111111110000000",
	"0000000000000000000000000000000000111111111111111111111100000000",
	"0000000000000000000000000000000001111111111111111111111000000000",
	"0000000000000000000000000000000011111111111111111111111000000000",
	"0000000000000000000000000000000111111111111111111111110000000000",
	"0000000000000000000000000000001111111111111111111111100000000000",
	"0000000000000000000000000000011111111111111111111111000000000000",
	"0000000000000000000000000000111111111111111111111110000000000000",
	"0000000000000000000000000001111111111111111111111110000000000000",
	"0000000000000000000000000011111111111111111111111100000000000000",
	"0000000000000000000000000111111111111111111111111000000000000000",
	"0000000000000000000000001111111111111111111111110000000000000000",
	"0000000000000000000000011111111111111111111111100000000000000000",
	"0000000000000000000000111111111111111111111111000000000000000000",
	"0000000000000000000001111111111111111111111110000000000000000000",
	"0000000000000000000011111111111111111111111000000000000000000000",
	"0000000000000000000111111111111111111111110000000000000000000000",
	"0000000000000000001111111111111111111111100000000000000000000000",
	"0000000000000000011111111111111111111111000000000000000000000000",
	"0000000000000000111111111111111111111110000000000000000000000000",
	"0000000000000001111111111111111111111100000000000000000000000000",
	"0000000000000001111111111111111111111000000000000000000000000000",
	"0000000000000011111111111111111111110000000000000000000000000000",
	"0000000000000111111111111111111111100000000000000000000000000000",
	"0000000000001111111111111111111111000000000000000000000000000000",
	"0000000000011111111111111111111110000000000000000000000000000000",
	"0000000000111111111111111111111100000000000000000000000000000000",
	"0000000000111111111111111111111000000000000000000000000000000000",
	"0000000001111111111111111111111000000000000000000000000000000000",
	"0000000011111111111111111111110000000000000000000000000000000000",
	"0000000011111111111111111111100000000000000000000000000000000000",
	"0000000111111111111111111111100000000000000000000000000000000000",
	"0000000111111111111111111111111111111111111111111111111111111110",
	"0000001111111111111111111111111111111111111111111111111111111110",
	"0000011111111111111111111111111111111111111111111111111111111110",
	"0000011111111111111111111111111111111111111111111111111111111110",
	"0000011111111111111111111111111111111111111111111111111111111110",
	"0000111111111111111111111111111111111111111111111111111111111110",
	"0000111111111111111111111111111111111111111111111111111111111110",
	"0001111111111111111111111111111111111111111111111111111111111110",
	"0001111111111111111111111111111111111111111111111111111111111110",
	"0001111111111111111111111111111111111111111111111111111111111110",
	"0011111111111111111111111111111111111111111111111111111111111110",
	"0011111111111111111111111111111111111111111111111111111111111110",
	"0011111111111111111111111111111111111111111111111111111111111110",
	"0011111111111111111111111111111111111111111111111111111111111110",
	"0011111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110",
	"0111111111111111111111111111111111111111111111111111111111111110");
	
	
	constant digito3 : digito := (
	"0000000000000000000000000011111111111100000000000000000000000000",
	"0000000000000000000001111111111111111111110000000000000000000000",
	"0000000000000000000111111111111111111111111100000000000000000000",
	"0000000000000000011111111111111111111111111111000000000000000000",
	"0000000000000001111111111111111111111111111111110000000000000000",
	"0000000000000011111111111111111111111111111111111000000000000000",
	"0000000000001111111111111111111111111111111111111100000000000000",
	"0000000000011111111111111111111111111111111111111110000000000000",
	"0000000000111111111111111111111111111111111111111111000000000000",
	"0000000001111111111111111111111111111111111111111111100000000000",
	"0000000001111111111111111111111111111111111111111111110000000000",
	"0000000011111111111111111111111111111111111111111111111000000000",
	"0000000111111111111111111111111111111111111111111111111000000000",
	"0000000111111111111111111111111111111111111111111111111100000000",
	"0000001111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111111111111111111111111111111110000000",
	"0000011111111111111111111111100000011111111111111111111110000000",
	"0000011111111111111111111110000000001111111111111111111111000000",
	"0000011111111111111111111100000000000011111111111111111111000000",
	"0000111111111111111111111000000000000011111111111111111111000000",
	"0000111111111111111111110000000000000001111111111111111111100000",
	"0000111111111111111111110000000000000001111111111111111111100000",
	"0000111111111111111111100000000000000000111111111111111111100000",
	"0001111111111111111111100000000000000000111111111111111111100000",
	"0001111111111111111111100000000000000000111111111111111111100000",
	"0000111111111111111111000000000000000000111111111111111111100000",
	"0000000000011111111111000000000000000000111111111111111111100000",
	"0000000000000000001111000000000000000000111111111111111111100000",
	"0000000000000000000000000000000000000000111111111111111111100000",
	"0000000000000000000000000000000000000000111111111111111111000000",
	"0000000000000000000000000000000000000001111111111111111111000000",
	"0000000000000000000000000000000000000001111111111111111111000000",
	"0000000000000000000000000000000000000001111111111111111110000000",
	"0000000000000000000000000000000000000011111111111111111110000000",
	"0000000000000000000000000000000000000111111111111111111100000000",
	"0000000000000000000000000000000000001111111111111111111100000000",
	"0000000000000000000000000000000000011111111111111111111000000000",
	"0000000000000000000000000000000011111111111111111111110000000000",
	"0000000000000000000000000000111111111111111111111111100000000000",
	"0000000000000000000000000001111111111111111111111111000000000000",
	"0000000000000000000000000001111111111111111111111110000000000000",
	"0000000000000000000000000001111111111111111111111100000000000000",
	"0000000000000000000000000001111111111111111111111000000000000000",
	"0000000000000000000000000001111111111111111111100000000000000000",
	"0000000000000000000000000001111111111111111110000000000000000000",
	"0000000000000000000000000001111111111111111111100000000000000000",
	"0000000000000000000000000001111111111111111111111100000000000000",
	"0000000000000000000000000001111111111111111111111111000000000000",
	"0000000000000000000000000001111111111111111111111111100000000000",
	"0000000000000000000000000011111111111111111111111111111000000000",
	"0000000000000000000000000011111111111111111111111111111100000000",
	"0000000000000000000000000011111111111111111111111111111110000000",
	"0000000000000000000000000011100000001111111111111111111111000000",
	"0000000000000000000000000000000000000011111111111111111111100000",
	"0000000000000000000000000000000000000000111111111111111111100000",
	"0000000000000000000000000000000000000000111111111111111111110000",
	"0000000000000000000000000000000000000000011111111111111111110000",
	"0000000000000000000000000000000000000000001111111111111111111000",
	"0000000000000000000000000000000000000000001111111111111111111000",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000000111111111111111111100",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000111100000000000000000000000011111111111111111110",
	"0000000111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111110000000000000000000000011111111111111111110",
	"0111111111111111111110000000000000000000000111111111111111111110",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111111000000000000000000000111111111111111111100",
	"0011111111111111111111000000000000000000001111111111111111111100",
	"0011111111111111111111100000000000000000001111111111111111111100",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111110000000000000000111111111111111111111000",
	"0001111111111111111111111000000000000001111111111111111111111000",
	"0000111111111111111111111110000000000011111111111111111111110000",
	"0000111111111111111111111111100000011111111111111111111111110000",
	"0000011111111111111111111111111111111111111111111111111111100000",
	"0000011111111111111111111111111111111111111111111111111111100000",
	"0000001111111111111111111111111111111111111111111111111111000000",
	"0000001111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000000001111111111111111111111111111111111111110000000000000",
	"0000000000000111111111111111111111111111111111111100000000000000",
	"0000000000000001111111111111111111111111111111110000000000000000",
	"0000000000000000011111111111111111111111111111100000000000000000",
	"0000000000000000000111111111111111111111111110000000000000000000",
	"0000000000000000000001111111111111111111110000000000000000000000",
	"0000000000000000000000000011111111111100000000000000000000000000");
	

	constant digito4 : digito := (
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000111111111111111100000000",
	"0000000000000000000000000000000000000001111111111111111100000000",
	"0000000000000000000000000000000000000001111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000111111111111111111100000000",
	"0000000000000000000000000000000000000111111111111111111100000000",
	"0000000000000000000000000000000000001111111111111111111100000000",
	"0000000000000000000000000000000000011111111111111111111100000000",
	"0000000000000000000000000000000000011111111111111111111100000000",
	"0000000000000000000000000000000000111111111111111111111100000000",
	"0000000000000000000000000000000001111111111111111111111100000000",
	"0000000000000000000000000000000001111111111111111111111100000000",
	"0000000000000000000000000000000011111111111111111111111100000000",
	"0000000000000000000000000000000111111111111111111111111100000000",
	"0000000000000000000000000000001111111111111111111111111100000000",
	"0000000000000000000000000000001111111111111111111111111100000000",
	"0000000000000000000000000000011111111111111111111111111100000000",
	"0000000000000000000000000000111111111111111111111111111100000000",
	"0000000000000000000000000000111111111111111111111111111100000000",
	"0000000000000000000000000001111111111111111111111111111100000000",
	"0000000000000000000000000011111111111111111111111111111100000000",
	"0000000000000000000000000011111111111111111111111111111100000000",
	"0000000000000000000000000111111111111111111111111111111100000000",
	"0000000000000000000000001111111111111111111111111111111100000000",
	"0000000000000000000000001111111111111111111111111111111100000000",
	"0000000000000000000000011111111111111111111111111111111100000000",
	"0000000000000000000000111111111111111111111111111111111100000000",
	"0000000000000000000000111111111111111111111111111111111100000000",
	"0000000000000000000001111111111111111111111111111111111100000000",
	"0000000000000000000011111111111111111011111111111111111100000000",
	"0000000000000000000011111111111111110011111111111111111100000000",
	"0000000000000000000111111111111111110011111111111111111100000000",
	"0000000000000000001111111111111111100011111111111111111100000000",
	"0000000000000000011111111111111111000011111111111111111100000000",
	"0000000000000000011111111111111111000011111111111111111100000000",
	"0000000000000000111111111111111110000011111111111111111100000000",
	"0000000000000001111111111111111100000011111111111111111100000000",
	"0000000000000001111111111111111000000011111111111111111100000000",
	"0000000000000011111111111111111000000011111111111111111100000000",
	"0000000000000111111111111111110000000011111111111111111100000000",
	"0000000000000111111111111111100000000011111111111111111100000000",
	"0000000000001111111111111111100000000011111111111111111100000000",
	"0000000000011111111111111111000000000011111111111111111100000000",
	"0000000000011111111111111110000000000011111111111111111100000000",
	"0000000000111111111111111110000000000011111111111111111100000000",
	"0000000001111111111111111100000000000011111111111111111100000000",
	"0000000001111111111111111000000000000011111111111111111100000000",
	"0000000011111111111111111000000000000011111111111111111100000000",
	"0000000111111111111111110000000000000011111111111111111100000000",
	"0000000111111111111111100000000000000011111111111111111100000000",
	"0000001111111111111111100000000000000011111111111111111100000000",
	"0000011111111111111111000000000000000011111111111111111100000000",
	"0000111111111111111110000000000000000011111111111111111100000000",
	"0000111111111111111110000000000000000011111111111111111100000000",
	"0001111111111111111100000000000000000011111111111111111100000000",
	"0011111111111111111000000000000000000011111111111111111100000000",
	"0011111111111111110000000000000000000011111111111111111100000000",
	"0111111111111111110000000000000000000011111111111111111100000000",
	"1111111111111111100000000000000000000011111111111111111100000000",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000011111111111111111100000000",
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000");
	
	
	constant digito5 : digito := (
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000111111111111111111111111111111111111111111111110000",
	"0000000000000111111111111111111111111111111111111111111111110000",
	"0000000000001111111111111111111111111111111111111111111111110000",
	"0000000000001111111111111111111111111111111111111111111111110000",
	"0000000000001111111111111111111111111111111111111111111111110000",
	"0000000000001111111111111111111111111111111111111111111111110000",
	"0000000000001111111111111111111111111111111111111111111111110000",
	"0000000000011111111111111111111111111111111111111111111111110000",
	"0000000000011111111111111111111111111111111111111111111111110000",
	"0000000000011111111111111111111111111111111111111111111111110000",
	"0000000000011111111111111111111111111111111111111111111111110000",
	"0000000000011111111111111111111111111111111111111111111111110000",
	"0000000000111111111111111111111111111111111111111111111111110000",
	"0000000000111111111111111111111111111111111111111111111111110000",
	"0000000000111111111111111111111111111111111111111111111111110000",
	"0000000000111111111111111111111111111111111111111111111111110000",
	"0000000000111111111111111111111111111111111111111111111111110000",
	"0000000001111111111111111111111111111111111111111111111111110000",
	"0000000001111111111111111111111111111111111111111111111111110000",
	"0000000001111111111111111111000000000000000000000000000000000000",
	"0000000001111111111111111111000000000000000000000000000000000000",
	"0000000001111111111111111111000000000000000000000000000000000000",
	"0000000011111111111111111110000000000000000000000000000000000000",
	"0000000011111111111111111110000000000000000000000000000000000000",
	"0000000011111111111111111110000000000000000000000000000000000000",
	"0000000011111111111111111110000000000000000000000000000000000000",
	"0000000111111111111111111110000000000000000000000000000000000000",
	"0000000111111111111111111100000000000000000000000000000000000000",
	"0000000111111111111111111100000000000000000000000000000000000000",
	"0000000111111111111111111100000000000000000000000000000000000000",
	"0000000111111111111111111100000000000000000000000000000000000000",
	"0000001111111111111111111000000000000000000000000000000000000000",
	"0000001111111111111111111000000011111111110000000000000000000000",
	"0000001111111111111111111000011111111111111110000000000000000000",
	"0000001111111111111111111011111111111111111111110000000000000000",
	"0000001111111111111111111111111111111111111111111100000000000000",
	"0000011111111111111111111111111111111111111111111110000000000000",
	"0000011111111111111111111111111111111111111111111111100000000000",
	"0000011111111111111111111111111111111111111111111111110000000000",
	"0000011111111111111111111111111111111111111111111111111000000000",
	"0000011111111111111111111111111111111111111111111111111100000000",
	"0000111111111111111111111111111111111111111111111111111110000000",
	"0000111111111111111111111111111111111111111111111111111111000000",
	"0000111111111111111111111111111111111111111111111111111111000000",
	"0000111111111111111111111111111111111111111111111111111111100000",
	"0000111111111111111111111111111111111111111111111111111111110000",
	"0001111111111111111111111111111111111111111111111111111111110000",
	"0001111111111111111111111111111111111111111111111111111111111000",
	"0001111111111111111111111111000000001111111111111111111111111000",
	"0001111111111111111111111000000000000011111111111111111111111100",
	"0011111111111111111111100000000000000000111111111111111111111100",
	"0011111111111111111111000000000000000000011111111111111111111100",
	"0011111111111111111110000000000000000000001111111111111111111110",
	"0000000111111111111100000000000000000000000111111111111111111110",
	"0000000000000001111000000000000000000000000111111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111110",
	"0000000000000000000000000000000000000000000011111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000000000000000000000000000000000000001111111111111111111",
	"0000000000001111000000000000000000000000000001111111111111111111",
	"0000111111111111000000000000000000000000000001111111111111111111",
	"1111111111111111000000000000000000000000000001111111111111111111",
	"1111111111111111100000000000000000000000000011111111111111111110",
	"1111111111111111100000000000000000000000000011111111111111111110",
	"0111111111111111110000000000000000000000000011111111111111111110",
	"0111111111111111110000000000000000000000000111111111111111111110",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000001111111111111111111100",
	"0011111111111111111100000000000000000000011111111111111111111100",
	"0011111111111111111110000000000000000000111111111111111111111000",
	"0011111111111111111111100000000000000001111111111111111111111000",
	"0001111111111111111111110000000000000111111111111111111111110000",
	"0001111111111111111111111110000000111111111111111111111111110000",
	"0000111111111111111111111111111111111111111111111111111111100000",
	"0000111111111111111111111111111111111111111111111111111111100000",
	"0000011111111111111111111111111111111111111111111111111111000000",
	"0000001111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111110000000000",
	"0000000000111111111111111111111111111111111111111111100000000000",
	"0000000000011111111111111111111111111111111111111111000000000000",
	"0000000000000111111111111111111111111111111111111100000000000000",
	"0000000000000011111111111111111111111111111111111000000000000000",
	"0000000000000000111111111111111111111111111111100000000000000000",
	"0000000000000000001111111111111111111111111110000000000000000000",
	"0000000000000000000001111111111111111111110000000000000000000000",
	"0000000000000000000000000111111111111100000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000");
	
	constant digito6 : digito := (
	"0000000000000000000000000000111111111110000000000000000000000000",
	"0000000000000000000000001111111111111111111000000000000000000000",
	"0000000000000000000001111111111111111111111111000000000000000000",
	"0000000000000000000111111111111111111111111111100000000000000000",
	"0000000000000000011111111111111111111111111111111000000000000000",
	"0000000000000000111111111111111111111111111111111100000000000000",
	"0000000000000011111111111111111111111111111111111110000000000000",
	"0000000000000111111111111111111111111111111111111111000000000000",
	"0000000000001111111111111111111111111111111111111111100000000000",
	"0000000000011111111111111111111111111111111111111111110000000000",
	"0000000000111111111111111111111111111111111111111111111000000000",
	"0000000000111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111000000011111111111111111111111000000",
	"0000001111111111111111111100000000001111111111111111111111000000",
	"0000011111111111111111111000000000000011111111111111111111100000",
	"0000011111111111111111110000000000000001111111111111111111100000",
	"0000111111111111111111100000000000000001111111111111111111100000",
	"0000111111111111111111000000000000000000111111111111111111100000",
	"0000111111111111111110000000000000000000111111111111111111110000",
	"0001111111111111111110000000000000000000111111111111111111110000",
	"0001111111111111111110000000000000000000011111111111111111110000",
	"0001111111111111111100000000000000000000011111111111111000000000",
	"0011111111111111111100000000000000000000011111000000000000000000",
	"0011111111111111111100000000000000000000000000000000000000000000",
	"0011111111111111111000000000000000000000000000000000000000000000",
	"0011111111111111111000000000000000000000000000000000000000000000",
	"0011111111111111111000000000000000000000000000000000000000000000",
	"0111111111111111111000000000000000000000000000000000000000000000",
	"0111111111111111111000000000000000000000000000000000000000000000",
	"0111111111111111110000000000000000000000000000000000000000000000",
	"0111111111111111110000000000000000000000000000000000000000000000",
	"0111111111111111110000000000001111111111000000000000000000000000",
	"0111111111111111110000000011111111111111111000000000000000000000",
	"0111111111111111110000001111111111111111111111000000000000000000",
	"1111111111111111110000011111111111111111111111110000000000000000",
	"1111111111111111110001111111111111111111111111111000000000000000",
	"1111111111111111110011111111111111111111111111111100000000000000",
	"1111111111111111110111111111111111111111111111111111000000000000",
	"1111111111111111111111111111111111111111111111111111100000000000",
	"1111111111111111111111111111111111111111111111111111110000000000",
	"1111111111111111111111111111111111111111111111111111111000000000",
	"1111111111111111111111111111111111111111111111111111111000000000",
	"1111111111111111111111111111111111111111111111111111111100000000",
	"1111111111111111111111111111111111111111111111111111111110000000",
	"1111111111111111111111111111111111111111111111111111111111000000",
	"1111111111111111111111111111111111111111111111111111111111000000",
	"1111111111111111111111111111111111111111111111111111111111100000",
	"1111111111111111111111111110000000111111111111111111111111100000",
	"1111111111111111111111111000000000000111111111111111111111110000",
	"1111111111111111111111110000000000000011111111111111111111110000",
	"1111111111111111111111100000000000000001111111111111111111110000",
	"1111111111111111111111000000000000000000111111111111111111111000",
	"1111111111111111111110000000000000000000011111111111111111111000",
	"1111111111111111111110000000000000000000011111111111111111111000",
	"1111111111111111111100000000000000000000001111111111111111111000",
	"1111111111111111111100000000000000000000001111111111111111111100",
	"1111111111111111111100000000000000000000001111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111000000000000000000000000111111111111111111100",
	"0011111111111111111000000000000000000000000111111111111111111100",
	"0011111111111111111000000000000000000000000111111111111111111100",
	"0011111111111111111000000000000000000000000111111111111111111100",
	"0011111111111111111100000000000000000000000111111111111111111100",
	"0011111111111111111100000000000000000000000111111111111111111100",
	"0001111111111111111100000000000000000000001111111111111111111000",
	"0001111111111111111110000000000000000000001111111111111111111000",
	"0001111111111111111110000000000000000000001111111111111111111000",
	"0000111111111111111111000000000000000000011111111111111111111000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111110000000000000000111111111111111111110000",
	"0000011111111111111111111000000000000001111111111111111111110000",
	"0000011111111111111111111100000000000111111111111111111111100000",
	"0000001111111111111111111111000000011111111111111111111111100000",
	"0000001111111111111111111111111111111111111111111111111111000000",
	"0000000111111111111111111111111111111111111111111111111111000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000011111111111111111111111111111111111111111111111110000000",
	"0000000001111111111111111111111111111111111111111111111100000000",
	"0000000000111111111111111111111111111111111111111111111000000000",
	"0000000000011111111111111111111111111111111111111111110000000000",
	"0000000000001111111111111111111111111111111111111111100000000000",
	"0000000000000111111111111111111111111111111111111111000000000000",
	"0000000000000011111111111111111111111111111111111110000000000000",
	"0000000000000001111111111111111111111111111111111100000000000000",
	"0000000000000000111111111111111111111111111111111000000000000000",
	"0000000000000000001111111111111111111111111111100000000000000000",
	"0000000000000000000011111111111111111111111110000000000000000000",
	"0000000000000000000000011111111111111111110000000000000000000000",
	"0000000000000000000000000011111111111100000000000000000000000000");
	
	
	constant digito7 : digito := (
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111100",
	"1111111111111111111111111111111111111111111111111111111111111000",
	"1111111111111111111111111111111111111111111111111111111111111000",
	"1111111111111111111111111111111111111111111111111111111111110000",
	"1111111111111111111111111111111111111111111111111111111111100000",
	"1111111111111111111111111111111111111111111111111111111111000000",
	"0000000000000000000000000000000000000000011111111111111110000000",
	"0000000000000000000000000000000000000000111111111111111100000000",
	"0000000000000000000000000000000000000001111111111111111000000000",
	"0000000000000000000000000000000000000011111111111111111000000000",
	"0000000000000000000000000000000000000011111111111111110000000000",
	"0000000000000000000000000000000000000111111111111111100000000000",
	"0000000000000000000000000000000000001111111111111111100000000000",
	"0000000000000000000000000000000000011111111111111111000000000000",
	"0000000000000000000000000000000000011111111111111110000000000000",
	"0000000000000000000000000000000000111111111111111110000000000000",
	"0000000000000000000000000000000001111111111111111100000000000000",
	"0000000000000000000000000000000001111111111111111000000000000000",
	"0000000000000000000000000000000011111111111111111000000000000000",
	"0000000000000000000000000000000111111111111111110000000000000000",
	"0000000000000000000000000000000111111111111111110000000000000000",
	"0000000000000000000000000000001111111111111111100000000000000000",
	"0000000000000000000000000000001111111111111111000000000000000000",
	"0000000000000000000000000000011111111111111111000000000000000000",
	"0000000000000000000000000000111111111111111110000000000000000000",
	"0000000000000000000000000000111111111111111110000000000000000000",
	"0000000000000000000000000001111111111111111100000000000000000000",
	"0000000000000000000000000001111111111111111100000000000000000000",
	"0000000000000000000000000011111111111111111000000000000000000000",
	"0000000000000000000000000011111111111111111000000000000000000000",
	"0000000000000000000000000111111111111111110000000000000000000000",
	"0000000000000000000000000111111111111111110000000000000000000000",
	"0000000000000000000000001111111111111111100000000000000000000000",
	"0000000000000000000000001111111111111111100000000000000000000000",
	"0000000000000000000000011111111111111111000000000000000000000000",
	"0000000000000000000000011111111111111111000000000000000000000000",
	"0000000000000000000000111111111111111111000000000000000000000000",
	"0000000000000000000000111111111111111110000000000000000000000000",
	"0000000000000000000000111111111111111110000000000000000000000000",
	"0000000000000000000001111111111111111100000000000000000000000000",
	"0000000000000000000001111111111111111100000000000000000000000000",
	"0000000000000000000011111111111111111100000000000000000000000000",
	"0000000000000000000011111111111111111000000000000000000000000000",
	"0000000000000000000011111111111111111000000000000000000000000000",
	"0000000000000000000111111111111111111000000000000000000000000000",
	"0000000000000000000111111111111111110000000000000000000000000000",
	"0000000000000000001111111111111111110000000000000000000000000000",
	"0000000000000000001111111111111111110000000000000000000000000000",
	"0000000000000000001111111111111111100000000000000000000000000000",
	"0000000000000000011111111111111111100000000000000000000000000000",
	"0000000000000000011111111111111111100000000000000000000000000000",
	"0000000000000000011111111111111111000000000000000000000000000000",
	"0000000000000000011111111111111111000000000000000000000000000000",
	"0000000000000000111111111111111111000000000000000000000000000000",
	"0000000000000000111111111111111111000000000000000000000000000000",
	"0000000000000000111111111111111110000000000000000000000000000000",
	"0000000000000001111111111111111110000000000000000000000000000000",
	"0000000000000001111111111111111110000000000000000000000000000000",
	"0000000000000001111111111111111110000000000000000000000000000000",
	"0000000000000001111111111111111100000000000000000000000000000000",
	"0000000000000001111111111111111100000000000000000000000000000000",
	"0000000000000011111111111111111100000000000000000000000000000000",
	"0000000000000011111111111111111100000000000000000000000000000000",
	"0000000000000011111111111111111100000000000000000000000000000000",
	"0000000000000011111111111111111100000000000000000000000000000000",
	"0000000000000011111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111111000000000000000000000000000000000",
	"0000000000000111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000001111111111111111110000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000",
	"0000000000000000000000000000000000000000000000000000000000000000");
	
	
	constant digito8 : digito := (
	"0000000000000000000000000111111111111110000000000000000000000000",
	"0000000000000000000011111111111111111111111000000000000000000000",
	"0000000000000000001111111111111111111111111111000000000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000011111111111111111111111111111111111100000000000000",
	"0000000000001111111111111111111111111111111111111111000000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111111111111111111111111111111111000000",
	"0000001111111111111111111111111111111111111111111111111111000000",
	"0000011111111111111111111111100000011111111111111111111111100000",
	"0000011111111111111111111110000000000111111111111111111111100000",
	"0000111111111111111111111000000000000001111111111111111111110000",
	"0000111111111111111111111000000000000000111111111111111111110000",
	"0000111111111111111111110000000000000000111111111111111111110000",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0000111111111111111111000000000000000000001111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0000011111111111111111100000000000000000011111111111111111100000",
	"0000011111111111111111110000000000000000111111111111111111100000",
	"0000011111111111111111110000000000000001111111111111111111000000",
	"0000001111111111111111111000000000000001111111111111111111000000",
	"0000000111111111111111111110000000000111111111111111111110000000",
	"0000000111111111111111111111100000011111111111111111111100000000",
	"0000000011111111111111111111111111111111111111111111111000000000",
	"0000000001111111111111111111111111111111111111111111110000000000",
	"0000000000111111111111111111111111111111111111111111100000000000",
	"0000000000001111111111111111111111111111111111111111000000000000",
	"0000000000000111111111111111111111111111111111111100000000000000",
	"0000000000000001111111111111111111111111111111111000000000000000",
	"0000000000000000001111111111111111111111111111000000000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000011111111111111111111111111111111111100000000000000",
	"0000000000001111111111111111111111111111111111111111000000000000",
	"0000000000011111111111111111111111111111111111111111100000000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000001111111111111111111111000000011111111111111111111111000000",
	"0000001111111111111111111100000000000011111111111111111111000000",
	"0000011111111111111111111000000000000001111111111111111111100000",
	"0000111111111111111111110000000000000000111111111111111111110000",
	"0000111111111111111111100000000000000000011111111111111111110000",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111000000000000000000001111111111111111111000",
	"0001111111111111111111000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111100000000000000000000000011111111111111111110",
	"0111111111111111111110000000000000000000000111111111111111111110",
	"0111111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111110000000000000000000000111111111111111111100",
	"0011111111111111111111000000000000000000000111111111111111111100",
	"0011111111111111111111000000000000000000001111111111111111111100",
	"0011111111111111111111100000000000000000001111111111111111111000",
	"0001111111111111111111100000000000000000011111111111111111111000",
	"0001111111111111111111110000000000000000111111111111111111111000",
	"0000111111111111111111111000000000000001111111111111111111110000",
	"0000111111111111111111111110000000000011111111111111111111110000",
	"0000011111111111111111111111100000001111111111111111111111100000",
	"0000011111111111111111111111111111111111111111111111111111100000",
	"0000001111111111111111111111111111111111111111111111111111000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000111111111111111111111111111111111111111111111111110000000",
	"0000000011111111111111111111111111111111111111111111111100000000",
	"0000000001111111111111111111111111111111111111111111111000000000",
	"0000000000111111111111111111111111111111111111111111110000000000",
	"0000000000001111111111111111111111111111111111111111100000000000",
	"0000000000000111111111111111111111111111111111111110000000000000",
	"0000000000000001111111111111111111111111111111111100000000000000",
	"0000000000000000111111111111111111111111111111110000000000000000",
	"0000000000000000000111111111111111111111111111000000000000000000",
	"0000000000000000000001111111111111111111111000000000000000000000",
	"0000000000000000000000000011111111111110000000000000000000000000");
	
	
	constant digito9 : digito := (
	"0000000000000000000000001111111111100000000000000000000000000000",
	"0000000000000000000011111111111111111110000000000000000000000000",
	"0000000000000000011111111111111111111111110000000000000000000000",
	"0000000000000001111111111111111111111111111100000000000000000000",
	"0000000000000011111111111111111111111111111111000000000000000000",
	"0000000000001111111111111111111111111111111111100000000000000000",
	"0000000000011111111111111111111111111111111111110000000000000000",
	"0000000000111111111111111111111111111111111111111000000000000000",
	"0000000001111111111111111111111111111111111111111100000000000000",
	"0000000011111111111111111111111111111111111111111110000000000000",
	"0000000111111111111111111111111111111111111111111111000000000000",
	"0000001111111111111111111111111111111111111111111111100000000000",
	"0000011111111111111111111111111111111111111111111111110000000000",
	"0000011111111111111111111111111111111111111111111111111000000000",
	"0000111111111111111111111111111111111111111111111111111000000000",
	"0000111111111111111111111111111111111111111111111111111100000000",
	"0001111111111111111111111110000001111111111111111111111100000000",
	"0001111111111111111111111000000000001111111111111111111110000000",
	"0011111111111111111111110000000000000111111111111111111110000000",
	"0011111111111111111111100000000000000011111111111111111111000000",
	"0011111111111111111111000000000000000001111111111111111111000000",
	"0111111111111111111110000000000000000000111111111111111111000000",
	"0111111111111111111110000000000000000000111111111111111111100000",
	"0111111111111111111100000000000000000000011111111111111111100000",
	"0111111111111111111100000000000000000000011111111111111111100000",
	"1111111111111111111100000000000000000000001111111111111111110000",
	"1111111111111111111000000000000000000000001111111111111111110000",
	"1111111111111111111000000000000000000000001111111111111111110000",
	"1111111111111111111000000000000000000000000111111111111111110000",
	"1111111111111111111000000000000000000000000111111111111111110000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111000",
	"1111111111111111111000000000000000000000000111111111111111111100",
	"1111111111111111111000000000000000000000000111111111111111111100",
	"0111111111111111111100000000000000000000000111111111111111111100",
	"0111111111111111111100000000000000000000001111111111111111111100",
	"0111111111111111111100000000000000000000001111111111111111111100",
	"0111111111111111111110000000000000000000001111111111111111111100",
	"0011111111111111111110000000000000000000011111111111111111111100",
	"0011111111111111111111000000000000000000011111111111111111111100",
	"0011111111111111111111000000000000000000111111111111111111111100",
	"0001111111111111111111100000000000000001111111111111111111111100",
	"0001111111111111111111110000000000000011111111111111111111111100",
	"0000111111111111111111111100000000000111111111111111111111111100",
	"0000111111111111111111111111000000111111111111111111111111111100",
	"0000011111111111111111111111111111111111111111111111111111111100",
	"0000001111111111111111111111111111111111111111111111111111111100",
	"0000001111111111111111111111111111111111111111111111111111111100",
	"0000000111111111111111111111111111111111111111111111111111111100",
	"0000000011111111111111111111111111111111111111111111111111111100",
	"0000000001111111111111111111111111111111111111111111111111111100",
	"0000000000111111111111111111111111111111111011111111111111111100",
	"0000000000001111111111111111111111111111110011111111111111111100",
	"0000000000000111111111111111111111111111100011111111111111111100",
	"0000000000000011111111111111111111111111000011111111111111111100",
	"0000000000000000111111111111111111111100000011111111111111111000",
	"0000000000000000000111111111111111110000000011111111111111111000",
	"0000000000000000000000111111111100000000000011111111111111111000",
	"0000000000000000000000000000000000000000000011111111111111111000",
	"0000000000000000000000000000000000000000000011111111111111111000",
	"0000000000000000000000000000000000000000000111111111111111111000",
	"0000000000000000000000000000000000000000000111111111111111111000",
	"0000000000000000000000000000000000000000000111111111111111110000",
	"0000000000000000000000000000000000000000000111111111111111110000",
	"0000000000000000000000000000000000000000000111111111111111110000",
	"0000000000000000000000000000000000000000001111111111111111110000",
	"0000000000000000111110000000000000000000001111111111111111110000",
	"0000000111111111111110000000000000000000001111111111111111100000",
	"0011111111111111111110000000000000000000011111111111111111100000",
	"0011111111111111111111000000000000000000011111111111111111100000",
	"0011111111111111111111000000000000000000011111111111111111000000",
	"0001111111111111111111000000000000000000111111111111111111000000",
	"0001111111111111111111100000000000000001111111111111111111000000",
	"0001111111111111111111100000000000000011111111111111111110000000",
	"0001111111111111111111110000000000000111111111111111111110000000",
	"0000111111111111111111111100000000001111111111111111111100000000",
	"0000111111111111111111111111000000111111111111111111111100000000",
	"0000111111111111111111111111111111111111111111111111111000000000",
	"0000011111111111111111111111111111111111111111111111111000000000",
	"0000011111111111111111111111111111111111111111111111110000000000",
	"0000001111111111111111111111111111111111111111111111100000000000",
	"0000001111111111111111111111111111111111111111111111000000000000",
	"0000000111111111111111111111111111111111111111111111000000000000",
	"0000000011111111111111111111111111111111111111111110000000000000",
	"0000000001111111111111111111111111111111111111111100000000000000",
	"0000000001111111111111111111111111111111111111111000000000000000",
	"0000000000111111111111111111111111111111111111100000000000000000",
	"0000000000011111111111111111111111111111111111000000000000000000",
	"0000000000000111111111111111111111111111111110000000000000000000",
	"0000000000000011111111111111111111111111111000000000000000000000",
	"0000000000000000111111111111111111111111100000000000000000000000",
	"0000000000000000001111111111111111111100000000000000000000000000",
	"0000000000000000000000111111111111000000000000000000000000000000");

	constant ponto1 : ponto :=(
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000001111111111111111111111111110000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000",
		"0000000000000000000000000000000000000000000000000000000000000000"
);	
-------------------------SINAIS DE CORES UTILIZADOS-------------------------------------------------	
signal color_red			: std_logic_vector (7 downto 0) :=("11100000");
constant color_white			: std_logic_vector (7 downto 0) :=("11111111");
-------------------------CONFIGURA��O 800 X 600-------------------------------------------------	
-------------------------CONFIGURA��O HORIZONTAL-------------------------------------------------	
constant h_area			: integer :=800;
constant h_frontporch	: integer :=40;
constant h_syncpulse		: integer :=128;
constant h_backporch		: integer :=88;
constant h_wholeline		: integer :=1056;
-------------------------CONFIGURA��O VERTICAL-------------------------------------------------
constant v_area				: integer :=600;
constant v_frontporch	: integer :=1;
constant v_syncpulse	: integer :=4;
constant v_backporch		: integer :=23;
constant v_wholeline		: integer :=628;
constant h_ajuste 		: integer:= 216;
constant v_ajuste 			: integer:= 27;

begin
	process (clk) 
-------------------------VARI�VEIS DE CONTAGEM-------------------------------------------------
	variable horizontal : integer :=0; 
	variable vertical   : integer :=0; 
-------------------------VARI�VEIS PARA MOSTRAR OS N�MEROS------------------------------------
	variable matriz_digitoq0 : digito; 
	variable matriz_digitoq1 : digito;	
	variable matriz_digitoq2 : digito;	
	variable matriz_digitoq3 : digito;	
	
begin
if rising_edge(clk) then
	if (horizontal >= h_syncpulse+h_backporch ) and (horizontal < h_syncpulse+h_backporch+h_area )
	and (vertical >= v_syncpulse+v_backporch )and (vertical < v_syncpulse+v_backporch+v_area )then
		if (estado < 8) then	
-------------------------MOSTRA NUMEROS Q0 Q1 Q2 Q3 EM POSI��ES DIFERENTES--------------------------------------------
-------------------------VARREDURA DE TODO O MONITOR NA RESOLU��O 800X600----------------------------------------------
			if ((vertical>=260+v_ajuste)and(vertical<=460+v_ajuste)and(horizontal>=200+h_ajuste)and(horizontal<=300+h_ajuste)) then
-------------------------ESCREVE DIGITO Q0---------------------------------------------------------------------------					
				if(matriz_digitoq0(vertical-(310+v_ajuste))(horizontal-(215+h_ajuste))='1') then 
						if (q0 = 0 and q1 < 2) then
						corestovga <= color_red;	
						else
						corestovga <= color_white;
						end if;
					else
						corestovga<="00000011"; --COR DO FUNDO GERAL DO BLOCO (PRETO)
					end if;
-------------------------ESCREVE DIGITO Q1---------------------------------------------------------------------------					 
			elsif ((vertical>=260+v_ajuste)and(vertical<=460+v_ajuste)and(horizontal>=320+h_ajuste)and(horizontal<=420+h_ajuste)) then
					if(matriz_digitoq1(vertical-(310+v_ajuste))(horizontal-(335+h_ajuste))='1') then
						if (q0 = 0 and q1 < 2) then
							corestovga <= color_red;	
						else
							corestovga <= color_white;
						end if;							
					else
						corestovga<="00000011"; --COR DO FUNDO GERAL DO BLOCO (PRETO)
					end if;
-------------------------ESCREVE DIGITO PONTO---------------------------------------------------------------------------	
			elsif ((vertical>=260+v_ajuste)and(vertical<=460+v_ajuste)and(horizontal>=440+h_ajuste)and(horizontal<=540+h_ajuste)) then
					if(ponto1(vertical-(310+v_ajuste))(horizontal-(455+h_ajuste))='1') then
						if (q0 = 0 and q1 < 2) then
							corestovga <= color_red;	
						else
							corestovga <= color_white;
						end if;	
					else
						corestovga<="00000011"; --COR DO FUNDO GERAL DO BLOCO (PRETO)
					end if;
-------------------------ESCREVE DIGITO Q2---------------------------------------------------------------------------						
			elsif ((vertical>=260+v_ajuste)and(vertical<=460+v_ajuste)and(horizontal>=560+h_ajuste)and(horizontal<=660+h_ajuste)) then
					if(matriz_digitoq2(vertical-(310+v_ajuste))(horizontal-(575+h_ajuste))='1') then
						if (q0 = 0 and q1 < 2) then
							corestovga <= color_red;	
						else
							corestovga <= color_white;
						end if;
					else
						corestovga<="00000011"; --COR DO FUNDO GERAL DO BLOCO (PRETO)
					end if;	
-------------------------ESCREVE DIGITO Q3---------------------------------------------------------------------------						
			elsif ((vertical>=260+v_ajuste)and(vertical<=460+v_ajuste)and(horizontal>=680+h_ajuste)and(horizontal<=780+h_ajuste)) then
				if(matriz_digitoq3(vertical-(310+v_ajuste))(horizontal-(695+h_ajuste))='1') then
					if (q0 = 0 and q1 < 2) then
								corestovga <= color_red;	
					else
								corestovga <= color_white;
					end if;
				else
					corestovga<="00000011"; --COR DO FUNDO GERAL DO BLOCO
				end if;				
			end if;	
			else
			corestovga<="00000011"; --COR DE FUNDO (PRETO)
		end if;	
	else
	corestovga<="00000011"; --COR DE FUNDO (PRETO)
	end if;
		
	-------------------------ATUALIZA��O DOS VALORES PARA VARREDURA DO MONITOR---------------------------------------------		
	if (horizontal > 0 )and (horizontal < h_syncpulse+1 )	then
		sync_h <= '0';
	else
		sync_h <= '1';
	end if;
		
	if (vertical > 0 ) and (vertical < v_syncpulse+1 )then
		sync_v <= '0';
	else
		sync_v <= '1';
	end if;
		
	horizontal := horizontal+1; 
		
if (horizontal=h_wholeline) then
		vertical := vertical+1; 
		horizontal := 0;
	end if;
		
	if (vertical=v_wholeline) then
		vertical := 0;
	end if;
end if;	

	case q0 is
		when 0 =>matriz_digitoq0:=digito0; 
		when 1 =>matriz_digitoq0:=digito1; 
		when 2 =>matriz_digitoq0:=digito2; 
		when 3 =>matriz_digitoq0:=digito3; 
		when 4 =>matriz_digitoq0:=digito4; 
		when 5 =>matriz_digitoq0:=digito5; 
		when 6 =>matriz_digitoq0:=digito6; 
		when 7 =>matriz_digitoq0:=digito7; 
		when 8 =>matriz_digitoq0:=digito8; 
		when 9 =>matriz_digitoq0:=digito9; 
		when others=>matriz_digitoq0:=digito0;  
	end case;

	case q1 is
		when 0 =>matriz_digitoq1:=digito0; 
		when 1 =>matriz_digitoq1:=digito1; 
		when 2 =>matriz_digitoq1:=digito2; 
		when 3 =>matriz_digitoq1:=digito3; 
		when 4 =>matriz_digitoq1:=digito4; 
		when 5 =>matriz_digitoq1:=digito5; 
		when 6 =>matriz_digitoq1:=digito6; 
		when 7 =>matriz_digitoq1:=digito7; 
		when 8 =>matriz_digitoq1:=digito8; 
		when 9 =>matriz_digitoq1:=digito9; 
		when others=>matriz_digitoq1:=digito0;  
	end case;

	case q2 is
		when 0 =>matriz_digitoq2:=digito0; 
		when 1 =>matriz_digitoq2:=digito1; 
		when 2 =>matriz_digitoq2:=digito2; 
		when 3 =>matriz_digitoq2:=digito3; 
		when 4 =>matriz_digitoq2:=digito4; 
		when 5 =>matriz_digitoq2:=digito5; 
		when others=>matriz_digitoq2:=digito0;  
	end case;

	case q3 is
		when 0 =>matriz_digitoq3:=digito0; 
		when 1 =>matriz_digitoq3:=digito1; 
		when 2 =>matriz_digitoq3:=digito2; 
		when 3 =>matriz_digitoq3:=digito3; 
		when 4 =>matriz_digitoq3:=digito4; 
		when 5 =>matriz_digitoq3:=digito5; 
		when 6 =>matriz_digitoq3:=digito6; 
		when 7 =>matriz_digitoq3:=digito7; 
		when 8 =>matriz_digitoq3:=digito8; 
		when 9 =>matriz_digitoq3:=digito9; 
		when others=>matriz_digitoq3:=digito0;  
	end case;
	

end process;


-------------------------PROCESSO PARA PISCAR NUMEROS QUANDO ESGOTA O TEMPO----------------------------	
process(clk1hz)
	variable cont: integer:=0;
begin
   if rising_edge(clk1hz) then
		if cont = 0 then    --CONT VARIANDO DE 0 PARA 1 A CADA PULSO DE CLOCK
		cont := cont+1;
		elsif cont > 0 then
			cont := 0;
      end if;
	end if; 
-------------------SE O TEMPO ESGOTAR O VALOR DE COLOR RED IRA MUDAR DE ACORDO COM CONT---------------------  
	if (q0 = 0 and q1 = 0 and q2 = 0 and q3 = 0) and flag_fim ='1' then
		if cont = 0 then
			color_red <= "11111111";
		elsif cont = 1 then
			color_red <= "11100000";
		end if;
	end if;		
end process;

end hardware;

